//================================================================
//     Custom String module
//		 
//		 This module is a submodule of Memory Management Module, it
//		 contains custom strings configurations to be displayed as  
//		 data chunks to screen
//================================================================
module Long_Strings(
	input VGA_CLK,
	input [4:0] String_Address,
	output reg[71:0] String_Data
);

always @(posedge VGA_CLK)
	begin
	case(String_Address)
	// Streaming
	00: String_Data <= 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
	01: String_Data <= 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
	02: String_Data <= 72'b011111000001000000000000000000000000000000000000001100000000000000000000;
	03: String_Data <= 72'b110001100011000000000000000000000000000000000000001100000000000000000000;
	04: String_Data <= 72'b110001100011000000000000000000000000000000000000000000000000000000000000;
	05: String_Data <= 72'b011000001111110011011100011111000111100011100110011100110111000111011000;
	06: String_Data <= 72'b001110000011000001110110110001100000110011111111001100011001101100110000;
	07: String_Data <= 72'b000011000011000001100110111111100111110011011011001100011001101100110000;
	08: String_Data <= 72'b000001100011000001100000110000001100110011011011001100011001101100110000;
	09: String_Data <= 72'b110001100011000001100000110000001100110011011011001100011001101100110000;
	10: String_Data <= 72'b110001100011011001100000110001101100110011011011001100011001101100110000;
	11: String_Data <= 72'b011111000001110011110000011111000111011011011011011110011001100111110000;
	12: String_Data <= 72'b000000000000000000000000000000000000000000000000000000000000000000110000;
	13: String_Data <= 72'b000000000000000000000000000000000000000000000000000000000000001100110000;
	14: String_Data <= 72'b000000000000000000000000000000000000000000000000000000000000000111100000;
	15: String_Data <= 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
	// Vp-p
	17: String_Data <= 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
	18: String_Data <= 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
	19: String_Data <= 72'b110000110000000000000000000000000000000000000000000000000000000000000000;
	20: String_Data <= 72'b110000110000000000000000000000000000000000000000000000000000000000000000;
	21: String_Data <= 72'b110000110000000000000000000000000000000000000000000000000000000000000000;
	22: String_Data <= 72'b110000110111110000000000011111000000000000000000000000000000000000000000;
	23: String_Data <= 72'b110000110110011000000000011001100000000000000000000000000000000000000000;
	24: String_Data <= 72'b110000110110011000000000011001100000000000000000000000000000000000000000;
	25: String_Data <= 72'b110000110110011000000000011001100000000000000000000000000000000000000000;
	26: String_Data <= 72'b011001100110011001111110011001100000000000000000000000000000000000000000;
	27: String_Data <= 72'b001111000110011000000000011001100000000000000000000000000000000000000000;
	28: String_Data <= 72'b000110000111110000000000011111000000000000000000000000000000000000000000;
	29: String_Data <= 72'b000000000110000000000000011000000000000000000000000000000000000000000000;
	30: String_Data <= 72'b000000000110000000000000011000000000000000000000000000000000000000000000;
	31: String_Data <= 72'b000000001111000000000000111100000000000000000000000000000000000000000000;
	32: String_Data <= 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase
	end
endmodule 